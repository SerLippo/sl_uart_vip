`ifndef UART_IF_SV
`define UART_IF_SV

interface uart_if;

  logic sdata;
  logic clk;

endinterface: uart_if

`endif