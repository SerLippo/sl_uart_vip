`ifndef UART_DEFINE_SV
`define UART_DEFINE_SV


`endif