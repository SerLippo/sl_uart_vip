`ifndef UART_TYPEDEF_SV
`define UART_TYPEDEF_SV

typedef enum {NONE, ODD, EVEN} uart_parity_kind_t;

`endif