`ifndef UART_TESTS_SVH
`define UART_TESTS_SVH

`include "uart_base_test.sv"
`include "uart_single_test.sv"
`include "uart_dual_test.sv"

`endif