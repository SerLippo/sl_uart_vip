`ifndef UART_SEQUENCES_SVH
`define UART_SEQUENCES_SVH

`include "uart_burst_seq.sv"

`include "uart_base_hseq.sv"
`include "uart_single_hseq.sv"


`endif